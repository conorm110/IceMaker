
);

endmodule
