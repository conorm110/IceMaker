
module REPLACE (
    